`timescale 1ms / 1ms

// Wrapper for interfacing with the MachXO2 Pico's hardware.
module machxo2_pico_frontend(
  // LEDs
  led0_n, // Pin M7/PB11A
  led1_n, // Pin N8/PB11B
  led2_n, // Pin B1/PL2A
  led3_n, // Pin B2/PL2B
  led4_n, // Pin C1/PL2C
  led5_n, // Pin C3/PL2D
  led6_n, // Pin C2/PL3A
  led7_n, // Pin D1/PL3B
  // Push-button
  button // Pin N3/PB6A
);

  // Clock frequency setup. Gives 0.992 Hz
  localparam OSCILLATOR_FREQ = "4.16"; // Oscillator freq, in MHz
  localparam FREQ_DIVIDER_BITS = 22; // Width of frequency divider counter

  input logic button;
  output logic led0_n, led1_n, led2_n, led3_n;
  output logic led4_n, led5_n, led6_n, led7_n;

  logic fast_clock; // approx 4.16 MHz, generated by internal oscillator
  logic slow_clock; // approx 0.992 Hz, generated from fast_clock by frequency divider
  logic reset_n;
  logic start;
  logic [3:0] multiplicand, multiplier;
  logic [7:0] product;

  // No reset button, so just keep it disabled.
  assign reset_n = 1'd1;

  // Multiplier inputs are hard-coded.
  assign multiplicand = 4'd11;
  assign multiplier = 4'd6;

  // LEDs show state of 'product'. They are active low.
  assign {led7_n, led6_n, led5_n, led4_n, led3_n, led2_n, led1_n, led0_n} = ~product;

  // Internal oscillator.
  OSCH #(.NOM_FREQ(OSCILLATOR_FREQ)) oscillator (
    .STDBY(1'd0),
    .OSC(fast_clock),
    .SEDSTDBY()
  );

  // Start button debouncer.
  debouncer start_debouncer (
    .clock(fast_clock),
    .reset_n(reset_n),
    .in(button),
    .out(start)
  );

  // Frequency divider to reduce fast 4.16 MHz clock to slow 0.992 Hz clock.
  freq_divider #(.BITS(FREQ_DIVIDER_BITS)) freq_divider (
    .in_clock(fast_clock),
    .out_clock(slow_clock),
    .reset_n(reset_n),
    .counter() // unused
  );

  // The actual 4-bit multiplier.
  multiplier #(.N(4)) mult (
    .clock(slow_clock),
    .reset_n(reset_n),
    .start(start),
    .ready(),
    .multiplicand(multiplicand),
    .multiplier(multiplier),
    .product(product)
  );
endmodule
