`timescale 1ms / 1ms

// Wrapper for interfacing with the MachXO2 Pico's hardware.
module machxo2_pico_frontend_8bit(
  // LEDs
  ledA0, // Pin M7/PB11A
  ledA1, // Pin N8/PB11B
  ledA2, // Pin B1/PL2A
  ledA3, // Pin B2/PL2B
  ledA4, // Pin C1/PL2C
  ledA5, // Pin C3/PL2D
  ledA6, // Pin C2/PL3A
  ledA7, // Pin D1/PL3B
  ledB0, // Pin N4/PB6D/SO
  ledB1, // Pin P13/PB20D/SI
  ledB2, // Pin P3/PB4C/CSS
  ledB3, // Pin B13/PT17C
  ledB4, // Pin A13/PT17D
  ledB5, // Pin C10/PT15D
  ledB6, // Pin K1/PL9A
  ledB7, // Pin K3/PL9B
  // Push-button
  button_n // Pin N3/PB6A
);

  // Clock frequency setup. Gives 0.992 Hz
  localparam OSCILLATOR_FREQ = "4.16"; // Oscillator freq, in MHz
  localparam FREQ_DIVIDER_BITS = 22; // Width of frequency divider counter
  localparam USE_SLOW_CLOCK = 1; // whether to use the slow clock instead of the fast clock for the multiplier

  input logic button_n;
  output logic ledA0, ledA1, ledA2, ledA3;
  output logic ledA4, ledA5, ledA6, ledA7;
  output logic ledB0, ledB1, ledB2, ledB3;
  output logic ledB4, ledB5, ledB6, ledB7;

  logic fast_clock; // approx 4.16 MHz, generated by internal oscillator
  logic slow_clock; // approx 0.992 Hz, generated from fast_clock by frequency divider
  logic reset_n;
  logic start, button;
  logic [7:0] multiplicand, multiplier;
  logic [15:0] product;

  // No reset button, so just keep it disabled.
  assign reset_n = 1'd1;

  assign button = ~button_n;

  // Multiplier inputs are hard-coded.
  assign multiplicand = 8'd45;
  assign multiplier = 8'd174;

  // LEDs show state of 'product'. They are active high.
  assign {ledA0, ledA1, ledA2, ledA3, ledA4, ledA5, ledA6, ledA7} = product[15:8];
  assign {ledB0, ledB1, ledB2, ledB3, ledB4, ledB5, ledB6, ledB7} = product[7:0];

  // Internal oscillator.
  OSCH #(.NOM_FREQ(OSCILLATOR_FREQ)) oscillator (
    .STDBY(1'd0),
    .OSC(fast_clock),
    .SEDSTDBY()
  );

  // Start button debouncer.
  debouncer start_debouncer (
    .clock(fast_clock),
    .reset_n(reset_n),
    .in(button),
    .out(start)
  );

  // Frequency divider to reduce fast 4.16 MHz clock to slow 0.992 Hz clock.
  freq_divider #(.BITS(FREQ_DIVIDER_BITS)) freq_divider (
    .in_clock(fast_clock),
    .out_clock(slow_clock),
    .reset_n(reset_n),
    .counter() // unused
  );

  // The actual 8-bit multiplier.
  multiplier #(.N(8)) mult (
    .clock(USE_SLOW_CLOCK ? slow_clock : fast_clock),
    .reset_n(reset_n),
    .start(start),
    .ready(),
    .multiplicand(multiplicand),
    .multiplier(multiplier),
    .product(product)
  );
endmodule
