`timescale 1ms / 1ms

// Wrapper for interfacing with the MachXO2 Pico's hardware.
module machxo2_pico_frontend(
  // LEDs
  led0, // Pin M7/PB11A
  led1, // Pin N8/PB11B
  led2, // Pin B1/PL2A
  led3, // Pin B2/PL2B
  led4, // Pin C1/PL2C
  led5, // Pin C3/PL2D
  led6, // Pin C2/PL3A
  led7, // Pin D1/PL3B
  // Push-button
  button_n // Pin N3/PB6A
);

  // Clock frequency setup. Gives 0.992 Hz
  localparam OSCILLATOR_FREQ = "4.16"; // Oscillator freq, in MHz
  localparam FREQ_DIVIDER_BITS = 22; // Width of frequency divider counter

  input logic button_n;
  output logic led0, led1, led2, led3;
  output logic led4, led5, led6, led7;

  logic fast_clock; // approx 4.16 MHz, generated by internal oscillator
  logic slow_clock; // approx 0.992 Hz, generated from fast_clock by frequency divider
  logic reset_n;
  logic start, ready, button;
  logic [3:0] multiplicand, multiplier;
  logic [7:0] product;

  // No reset button, so just keep it disabled.
  assign reset_n = 1'd1;

  assign button = ~button_n;

  // Multiplier inputs are hard-coded.
  assign multiplicand = 4'd11;
  assign multiplier = 4'd6;

  // LEDs show state of 'product'. They are active low.
  //assign {led0, led1, led2, led3, led4, led5, led6, led7} = product;
  assign {led0, led1, led2, led3, led4, led5, led6, led7} = {fast_clock, slow_clock, reset_n, button, start, ready, 1'd0};

  // Internal oscillator.
  OSCH #(.NOM_FREQ(OSCILLATOR_FREQ)) oscillator (
    .STDBY(1'd0),
    .OSC(fast_clock),
    .SEDSTDBY()
  );

  // Start button debouncer.
  debouncer start_debouncer (
    .clock(fast_clock),
    .reset_n(reset_n),
    .in(button),
    .out(start)
  );

  // Frequency divider to reduce fast 4.16 MHz clock to slow 0.992 Hz clock.
  freq_divider #(.BITS(FREQ_DIVIDER_BITS)) freq_divider (
    .in_clock(fast_clock),
    .out_clock(slow_clock),
    .reset_n(reset_n),
    .counter() // unused
  );

  // The actual 4-bit multiplier.
  multiplier #(.N(4)) mult (
    .clock(slow_clock),
    .reset_n(reset_n),
    .start(start),
    .ready(ready),
    .multiplicand(multiplicand),
    .multiplier(multiplier),
    .product(product)
  );
endmodule
